module prom_hd(addr,data_out);
input [15:0]addr;
output [26:0]data_out;
parameter mem_depth = 1 <<16; 

reg [26:0]prom_reg[65535:0];

initial
begin
								//$readmemb("rom_code_full",prom_reg);
								$display($time,"Starting HD with HD instruction");
								prom_reg[0] =  27'b1_0001_000_101_1000000000001011; //IMM ADD 
								prom_reg[1] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[2] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[3] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[4] =  27'b1_0001_001_101_0000000000001111; //IMM ADD
								prom_reg[5] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[6] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[7] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[8] =  27'b0_1011_010_000_0000000000000001; // reg HD
								prom_reg[9] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[10] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[11] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[12] =  27'b0_0000_000_000_0000000000000000; //NOP
								$display($time,"Done HD with HD instruction");
								$display($time,"Starting HD without HD instruction");
								prom_reg[13] =  27'b1_0001_000_101_1000000000001011; //IMM ADD (0) = A 
								prom_reg[14] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[15] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[16] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[17] =  27'b1_0001_001_101_0000000000001111; //IMM ADD  (1) = B
								prom_reg[18] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[19] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[20] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[21] =  27'b1_0001_010_101_0000000000000000; //IMM ADD (2) = 0
								prom_reg[22] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[23] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[24] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[25] =  27'b1_0001_011_101_0000000000010000; //IMM ADD (3) = 16
								prom_reg[26] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[27] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[28] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[29] =  27'b1_0001_100_101_0000000000000000; //IMM ADD (4) = 0
								prom_reg[30] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[31] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[32] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[33] =  27'b1_0110_101_000_0000000000000001; //IMM AND (5) = (0) & 1
								prom_reg[34] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[35] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[36] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[37] =  27'b1_0110_110_001_0000000000000001; //IMM AND (6) = (1) & 1
								prom_reg[38] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[39] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[40] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[41] =  27'b0_0001_111_101_0000000000000110; //REG ADD (7) = (5) + (6)
								prom_reg[42] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[43] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[44] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[45] =  27'b1_0110_111_111_0000000000000001; //IMM AND (7) = (7) & 1
								prom_reg[46] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[47] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[48] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[49] =  27'b0_0001_010_010_0000000000000111; //reg ADD (2) = (2) + (7)
								prom_reg[50] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[51] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[52] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[53] =  27'b1_0101_000_000_0000000000000001; //IMM LSR (0) = (0) >> 1 
								prom_reg[54] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[55] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[56] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[57] =  27'b1_0101_001_001_0000000000000001; //IMM LSR (1) = (1) >> 1 
								prom_reg[58] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[59] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[60] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[61] =  27'b1_0010_011_011_0000000000000001; //IMM SUB (3) = (3) -1
								prom_reg[62] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[63] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[64] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[65] =  27'b0_1101_011_100_1111111111101111; //BNEQ (3) (4) 
								prom_reg[66] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[67] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[68] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[69] =  27'b1_0000_000_000_0000000000000000; //HALT
								$display($time,"Done HD without HD instruction");
end         
assign data_out = prom_reg[addr];

endmodule
