module prom(addr,data_out);
input [15:0]addr;
output [26:0]data_out;
parameter mem_depth = 1 <<16; 

reg [26:0]prom_reg[65535:0];

initial
begin
								//$readmemb("rom_code_full",prom_reg);
								prom_reg[0] =  27'b1_0001_000_101_1111111111111111; //IMM ADD 
								prom_reg[1] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[2] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[3] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[4] =  27'b1_0001_001_000_0000000000001111; //IMM ADD
								prom_reg[5] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[6] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[7] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[8] =  27'b0_0001_010_000_0000000000000001; //REG ADD
								prom_reg[9] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[10] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[11] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[12] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[13] =  27'b1_0010_001_101_0000000000001110; //IMM SUB
								prom_reg[14] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[15] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[16] =  27'b0_0000_000_000_0000000000000000; //NOP 
								prom_reg[17] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[18] =  27'b0_0010_100_010_0000000000000001; // REG SUB 
								prom_reg[19] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[20] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[21] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[22] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[23] =  27'b1_0001_011_101_1000000000001010; //IMM ADD 
								prom_reg[24] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[25] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[26] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[27] =  27'b0_0011_110_011_0000000000000001; //reg ASR
								prom_reg[28] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[29] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[30] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[31] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[32] =  27'b1_0011_111_010_0000000000000011; //IMM ASR
								prom_reg[33] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[34] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[35] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[36] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[37] =  27'b0_0100_101_000_0000000000000111; //REG LSL
								prom_reg[38] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[39] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[40] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[41] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[42] =  27'b1_0100_111_010_0000000000000011; //IMM LSL
								prom_reg[43] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[44] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[45] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[46] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[47] =  27'b0_0101_000_011_0000000000000000; //REG LSR
								prom_reg[48] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[49] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[50] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[51] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[52] =  27'b1_0101_101_111_0000000000000001; //IMM LSR
								prom_reg[53] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[54] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[55] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[56] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[57] =  27'b0_0110_110_001_0000000000000010; //REG AND
								prom_reg[58] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[59] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[60] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[61] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[62] =  27'b1_0110_100_001_0000000001011001; //IMM AND
								prom_reg[63] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[64] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[65] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[66] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[67] =  27'b0_0111_111_010_0000000000000101; //REG OR
								prom_reg[68] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[69] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[70] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[71] =  27'b1_0111_010_000_0000000000000011; //IMM OR
								prom_reg[72] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[73] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[74] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[75] =  27'b0_1000_000_001_0000000000000010; //REG SLT
								prom_reg[76] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[77] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[78] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[79] =  27'b1_1000_000_001_0000000000001111; //IMM SLT
								prom_reg[80] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[81] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[82] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[83] =  27'b0_1001_001_000_0000000000000111; //    INV
								prom_reg[84] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[85] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[86] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[87] =  27'b1_1010_110_001_0000000000000111; // reg MOV
								prom_reg[88] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[89] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[90] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[91] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[92] =  27'b0_1010_111_000_0000000000011111; // IMM MOV
								prom_reg[93] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[94] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[95] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[96] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[97] =  27'b1_1011_010_010_0000000000000101; // reg HD
								prom_reg[98] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[99] =  27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[100] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[101] = 27'b0_1011_010_111_0000000000000111; // IMM HD
								prom_reg[102] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[103] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[104] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[105] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[106] = 27'b1_1111_01_001_00000000000000000; //	STORE BYTE
								prom_reg[107] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[108] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[109] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[110] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[111] = 27'b1_1111_00_101_00000000000000000; //	LOAD BYTE
								prom_reg[112] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[113] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[114] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[115] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[116] = 27'b1_1111_01_110_01000000000000001; //	STORE word
								prom_reg[117] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[118] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[119] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[120] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[121] = 27'b1_1111_10_100_00000000000000001; //	LOAD_WORD 
								prom_reg[122] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[123] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[124] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[125] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[126] = 27'b0_1100_111_111_0000000000000010; // BEQ
								prom_reg[127] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[128] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[129] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[130] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[131] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[132] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[133] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[134] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[135] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[136] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[137] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[138] = 27'b0_1100_111_110_0000000000000010; // BEQ
								prom_reg[139] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[140] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[141] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[142] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[143] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[144] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[145] = 27'b0_1101_101_111_0000000000000010; // BNEQ
								prom_reg[146] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[147] = 27'b0_0000_000_000_0000000000000000; //NOP
				 				prom_reg[148] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[149] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[150] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[151] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[152] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[153] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[154] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[155] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[156] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[157] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[158] = 27'b0_1110_000_000_0000000001010011; //jump
								prom_reg[159] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[160] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[161] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[162] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[163] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[164] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[165] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[166] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[167] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[168] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[169] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[170] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[171] = 27'b0_0000_000_000_0000000000000000; //NOP
								prom_reg[172] = 27'b1_0000_000_000_0000000000000000; //NOP
end         
assign data_out = prom_reg[addr];

endmodule
